module alu(
           input [3:0] A,B,  // ALU 4-bit Inputs
           input [3:0] ALU_Sel,// ALU Selection
           output [7:0] ALU_Out, // ALU 8-bit Output
           output CarryOut // Carry Out Flag
    );
    reg [7:0] ALU_Result;
    wire [8:0] tmp;
    assign ALU_Out = ALU_Result; // ALU out
    assign tmp = {1'b0,A} + {1'b0,B};
    assign CarryOut = tmp[8]; // Carryout flag
    always @(*)
    begin
        case(ALU_Sel)
        4'b0000: // Addition
           ALU_Result = A + B ;
        4'b0001: // Subtraction
           ALU_Result = A - B ;
        4'b0010: // Multiplication
           ALU_Result = A * B;
        4'b0011: // Division
           ALU_Result = A/B;
        4'b0100: // Logical shift left
           ALU_Result = A<<1;
         4'b0101: // Logical shift right
           ALU_Result = A>>1;
         4'b0110: // Rotate left
           ALU_Result = {A[6:0],A[7]};
         4'b0111: // Rotate right
           ALU_Result = {A[0],A[7:1]};
          4'b1000: //  Logical and
           ALU_Result = A & B;
          4'b1001: //  Logical or
           ALU_Result = A | B;
          4'b1010: //  Logical xor
           ALU_Result = A ^ B;
          4'b1011: //  Logical nor
           ALU_Result = ~(A | B);
          4'b1100: // Logical nand
           ALU_Result = ~(A & B);
          4'b1101: // Logical xnor
           ALU_Result = ~(A ^ B);
          4'b1110: // Greater comparison
           ALU_Result = (A>B)?8'd1:8'd0 ;
          4'b1111: // Equal comparison
            ALU_Result = (A==B)?8'd1:8'd0 ;
          default: ALU_Result = 0 ;
        endcase
    end

endmodule

//---------------------------------------------------------------
module TriBuff(en, rst, In, Ou);
input wire en;
input wire rst;
input wire [3:0] In;
output reg [3:0]Ou;

    if (rst == 1) begin
      Ou <= 0;
    end else if (rst == 0) begin
      if (en == 0) begin
        Ou <= 4'bzzzz;
      end else if (en == 1) begin
        Ou <= In;
      end
    end


endmodule
//-------------------------------------------------------------------
module accum (en, rst, In, Ou);
input wire rst;
input wire [3:0] In;
output reg [3:0]Ou;
reg [3:0] Ac;
Initial Ac <= 0;
if (rst == 0) begin
  Ou <= In + Ac;
end else begin
  Ou <=4'b0;
end
